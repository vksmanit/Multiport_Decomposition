*********** MP2 ***********
******* node 8 is gnd *******
R10 5 6 1k
I11 5 7 DC 1m
R12 6 0 1k
R13 7 0 1k
V1 5 6 DC 0
V2 6 7 DC 0
.end
