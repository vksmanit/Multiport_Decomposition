*************** ckt-04 *************
R1 1 2  2k
R2 1 3  2k
R3 2 3  2k
R4 2 4  2k
I5 3 4  DC 2m
R6 1 5  2k
R7 2 6  2k
R8 4 10 2k
R9 3 9  2k


R10 5 6 1k
I11 5 7 DC 1m
R12 6 8 1k
R13 7 8 1k


R14 9 10 3k
R15 9 11  3k
R16 10 11 3k
I17 11 13 DC 3m

R18 7 12  4k
R19 12 13 4k
R20 12 0  4k
R21 13 0  4k

.op
.control 
run 
*print all
print (v(1) - v(2))
print (v(1) - v(3))
print (v(2) - v(3))
print (v(2) - v(4))
print (v(3) - v(4))
print (v(1) - v(5))
print (v(2) - v(6))
print (v(4) - v(10))
print (v(3) - v(9))

print (v(5) - v(6))
print (v(5) - v(7))
print (v(6) - v(8))
print (v(7) - v(8))


print (v(9) - v(10))
print (v(9) - v(11))
print (v(10)- v(11))
print (v(11)- v(13))
print (v(7) - v(12))
print (v(12) - v(13))
print (v(12))
print (v(13))

.endc
.end
