*********** MP1 ************
***** node 10 is gnd *****88
R1 1 2  2k
R2 1 3  2k
R3 2 3  2k
R4 2 4  2k
I5 3 4  DC 2m
R6 1 5  2k
R7 2 6  2k
R8 4 0 2k
R9 3 9  2k
V1 5 6 DC 0
V2 6 9 DC 0
V3 9 0 DC 0
.end

