*****************888
r6 1 5 2k 
r7 3 6 2k 
r8 4 0 2k 
r9 5 6 2k 
r10 5 7 2k 
r11 6 7 2k 
r12 6 0 2k 
r13 7 0 2k
v1 1 3 DC 0
v2 3 4 DC 1
