R1 1 2  2k
R2 1 3  2k
R3 2 3  2k
R4 2 4  2k
I5 3 4  DC 2m
R6 1 5  2k
R7 2 6  2k
R8 4 0 2k
R9 3 9  2k


R10 5 6 1k
I11 5 7 DC 1m
R12 6 0 1k
R13 7 0 1k


R14 9 10 3k
R15 9 0  3k
R16 10 0 3k
I17 0 7 DC 3m

.control 
.op 
run 
print all
.endc
.end
