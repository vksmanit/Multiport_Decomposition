******* MP3 ************
****** node gnd is gnd ****
R14 9 10 3k
R15 9 0  3k
R16 10 0 3k
I17 0 7 DC 3m
V1 7 9 DC 0
V2 9 10 DC 0
.end
