*******************
i1 1 2 DC 1m
r2 1 3 1k 
r3 2 3 1k 
r4 2 4 1k 
r5 3 4 1k 
***********
r6  1 5 2k 
r7  4 0 2k 
r8  5 6 2k 
r9  5 7 2k 
r10 6 7 2k 
r11 6 0 2k 
r12 7 0 2k

.op 
.control
run 
print (v(1) - v(2))
print (v(1) - v(3))
print (v(2) - v(3))
print (v(2) - v(4))
print (v(3) - v(4))


print (v(1) - v(5))
print (v(4)       )
print (v(5) - v(6))
print (v(5) - v(7))
print (v(6) - v(7))
print (v(6)       )
print (v(7)       )

.endc
.end
